LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY HALFADDER IS
	PORT (
		A : IN STD_LOGIC;
		B : IN STD_LOGIC;
		SI : OUT STD_LOGIC;
		CI : OUT STD_LOGIC);
END HALFADDER;

ARCHITECTURE ARHA OF HALFADDER IS
BEGIN
	SI <= A XOR B;
	CI <= A AND B;
END ARHA;